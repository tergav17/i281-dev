������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: CAT FILE1 FILE2 ...
 CAN'T OPEN FILE
                                                               0 ��� �<^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��G4 �F0 ��� P ��48��;                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�0����0���0���0��0����r�l��48��pP �0�l0048��h0�l0 �48��aP �&0 4����� P �4 ��4����� � � ��4����0��0���0�����P��0 T8� �߀P��4 ���P�� � ��4 �0                                                                                      