������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
                                                                          0 ��� �<^8�8 �r�l��� 4 � �X��� P �0� �X��4-� �X� P �%4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��B4 �A0 ��� P ��0 �+48��44 �5�.48��.                                                                                        ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
 UNEXPECTED CHAR IN NUM
                                                                                      8�8�� 48��{8�8�� 48��t�P ��48��n                                                                                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�����r��� 4 ��4 � �48��t�P��0:48��m�,��-�8�� �0:48��b0 48��^�.p�@ P48��� �8 ���l48��N|8 �0'48��04�8��0 4d8��0 4
8��00�0 48��\�4������m �x�h ����< � �80�X����P ���48���                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0��0��|0 ���,�-0��0��P�� � ��r�l�8�8�48��dP �0�48��\4�l0 48��XP ��\�S|�� � �'��P ���� 4 ��P��X �8
��0 T�8� ��P��8�48��0P �0 4���\��0 �\�#                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8��P���-P�-��,P�,�P �h�<4
� �4���a�4;� �2X �4 � �-40� �49� �4��*4a� �4z� �p 4A� �4Z� �4���� �8 ��;X �94;� ���	4'� �4"� ��-��+8�� 48��/�8 � �8ܻ 48��&��40� �49� �4a� �4z� �p 4A� �4Z� �X4*� ����0 ��4���\�    