������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: DEBUG FILE
 CAN'T CREATE FILE
 OUT OF SPACE
 BAD RECORD
 
?
*                                   0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ��� p��8Ȼ 48��:48��7                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0W�0Z8�4�l48��z4�l48��u0 ���	8�� 48��jP ��4���4 ��X ��pQ48��\��0 ���4��� 4 ��X�40� �N49� �4A� �H4F� �Epp0���0E �J �Tp���H ��0���0��/                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 �8 4��� 4��� X�����r�l�8�48��pP �48��kP �0'�(0�l8 �
" 48��_P ��
0J4��� t��t���4@ �T� ��� T��4�� X��0��048��=4�4�l48��8                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |��4 ��4@ �T� ��� X �t��� 8 ���8�8�l48��iP �.4 ���4���0� 0��04�� P��4��0 8 � P��4	��0 8 � P��4
��0 � P���0;T �	�
�P�
�0��\�64 ��4�4�l48��.                                                                                    