������������������������������������������������������������������������������������������������������������������������������
 UA NAME   EX SIZE
 0:  *.*  FILES OVER   BLOCKS
 NO FILES
                                                                0 ��<^48�8��{48��v4
8��uP 0648��p0 ����	048��g�P���P��j4���4 ��048��V0�0 � �`48��N� �P� ���p�0.48��B0�0��0 48��:�	�iA �	��P�hA �0 8ٻ 48��(0 48��&48��#P ��48��4 �                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8 �P �0'48��04�8��0 4d8��
0 4
8��0 48��\�g�����h�im �x�h ��h�i�< � �80�X����P ���H48���F8�0 48��@��h��i08˻ ��048��4��h�	�i08׻ ��0,48��(4 �'                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �r�l��8 � 4 � �X��� P �� �X��04��p:�
�p �0*��0.�0 �" 48��\8 ���l48��V                                                                                                                                                                          