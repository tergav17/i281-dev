������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
 CAN'T OPEN FILE
                                                           0 ��� �<^8�8 �r�l��� 4 � �X��� P �.� �X��4-� �X� P �#4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��D4 �C0 ��� P ��0 �%48��64 �74���                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8�� 48��{8�8�� 48��t�P ��48��n                                                                                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0��0��|0 ���0��P�� � ��r�l�8�8�48��gP �0�l0448��]4�l0 48��YP ��\�T|�� � �'��P ���� 4 ��P��X �8
��0 T�8� ��P��8�48��1P �0 4���\��0 �\�$                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8��P �h�<4
� �4 ��a�4;� �2X �4 � �-40� �49� �4��*4a� �4z� �p 4A� �4Z� �4���� �8 ��;X �94;� ���	4'� �4"� ��-��+8�� 48��:�8� �8ѻ 48��1��40� �49� �4a� �4z� �p 4A� �4Z� �X4$� ����0 ��4���\�                          