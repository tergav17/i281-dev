������������������������������������������������������������������������������������������������������������������������������?:*.*  FILES IN USE
  BLOCKS IN USE
  BLOCKS FREE
                                                                           0 ��<^48�8��|0 ����	0�l0 4
8��qP ��P���P��	�iA �	��P�hA ��	P�	��P�48��T�� ��08�� 48��H048��F�� �	�08Ȼ 48��:048��848��5�n� �o�08ٻ 48��)0'48��'4 �&                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8 �P �0'48��04�8��0 4d8��0 4
8��00�0 48��\�f����� �m �x�h �� ��< � �80�X����P ���F48���E                                                                                                                                  