������������������������������������������������������������������������������������������������������������������������������
 UA NAME   EX SIZE
 0:  *.*  FILES OVER   BLOCKS
 NO FILES
                                                                0 ��<^48�8��|48��w4
8��v4�lP 0648��o0 ����	048��f�P���P��j4���4 ��048��U0�0 � �`48��M� �P� ���p�0.48��A0�0��0 48��9�	�iA �	��P�hA �0 8ۻ 48��'0 48��%48��"P ��48��4 �                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8 �P �0'48��04�8��0 4d8��0 4
8��00�0 48��\�f�����h�im �x�h ��h�i�< � �80�X����P ���F48���E8�0 48��?��h��i08ͻ ��048��3��h�	�i08ٻ ��0,48��'4 �&                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �r�l��8 � 4 � �X��� P �� �X��04��p:�
�p �0*��0.�0 �" 48 ��8��[8 ���l48��U                                                                                                                                                                      