������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
  /FY 4                                                            0 ��� �<^8�8 �r�l��� 4 � �X��� P �0� �X��4-� �X� P �%4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��B4 �A0 ��� P ��0 �E48��44 �54 ���48��,                                                                                    ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
 UNEXPECTED CHAR IN NUMERIC
 UNDEFINED EXPRESSION
 UNEXPECTED TOKEN
 VALUE STACK OVERFLOW
                 8�8�� 48��{8�8�� 48��t�0P �
p���8�� 48��j����48��d                                                                                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������EXPRESSION STACK OVERFLOW
 VALUE STACK DEPLETION
 EXPRESSION STACK DEPLETION
                                                8��H��9�r��� 4 ��4 � �48��t�9P��0:48��m�F��G�8�� �0:48��b0 48��^�p�@ P48��� �8 ���l48��N|8 �0'48��04�8��0 4d8��0 4
8��00�0 48��\�4������m �x�h ����< � �80�X����P ���48���                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |4�8��5P�{�58��x0��10��60��5|0 �4�2�7�80�3�1P�1� � ��r�l�8�8�48��]P �	�1�H0 �F�G0�48��P4�l0 48��LP ��\�G|�1� � �'�4�3P ���� 4 ��P�4�6X �8
�6�0 T�38� ��2P��28�48��$P �0 4�3��\��0 �6\�                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �1�H�8P�8�7�T�7�F�G�6P �l�=4
� �4��5�e�54;� �3X �4 � �.40� �49� 4��,4a� �4z� �p 4_� �4A� �4Z� 4���5� �8 �5�>X �<4;� ��5�	4'� �4"� ��0�5�.8�� 48��1�08:� �98ڻ 48��(�9�640� �49� �4a� �4z� �p 4_� �4A� �4Z� �X4D� ����0 ��4��6�0\�  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0
�0 ��0:� T �wt0�	4�P� 89� �P�( � T �X����t9�T9�90 ���98tX�t��
8t�8t��0�48��N��9� P �J����|�	�B ���PA �����9� P40� ��49� �4A� ��4F� ��xx0�� �ӄF ��ԄT���                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0$�/0�.8��0p���<P �	�;pF�p��0 ���8�� 48��gp��0 ���p��0 ���/0)� 0���� ��T�/�p����.0� 0���0� ��T�.�0�48��=8�8̻ 48��6�0�p���p���p���p���48��)                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8p�)p�'8p��$p�"p�� 8pW�8p��8p��8p=�p�� p�p��"8�� 48��]�0�� 8�0�48��T��.4� �	���� �8�� 4	8��F48��C48��@0 \�>                                                                                                                      �	�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0��.8� �6t�.0��/8&� �/������������t�/�.� p+���A ����PA ��p���a ����pa ��p�� �/������\�G48��C                                                                                                                                  