������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: CP SOURCE DEST
                                                                                      0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ��� p��r�l�48��;P �0�l0 48��3�48��/P �0�l048��'0 ��0��48��                                                      ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN SOURCE FILE
 CAN'T CREATE DEST FILE
 CAN'T OPEN DEST FILE
 DEST WRITE ERROR
                                     8��r�l�48��|P �0 �?0 �@ @ P�l�48��nP �0 ��
�P����P�4 � ��r�l�48��YP �02�0 ��� �@ @ P�l�4	8��HP �0I��P��P���P ���4�l48��448��/                                                                                          