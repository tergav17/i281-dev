������������������������������������������������������������������������������������������������������������������������������NO ARGUMENT
 CAN'T OPEN FILE
                                                                                                 0 ��<^8��r�l��8 � 4 � �X��� P �� �
X��0 ��0�l0 48��e0 ��" 48��_P �0�l048��W0�l0 � 48��PP �0 4����� P �4 ��48��A��P��0 T8� �� P��4 �4                                                                                                