������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: XMODEM [-ST] FILE
 CAN'T OPEN FILE
 CAN'T CREATE FILE
 TRANSFER FAILED
                        0 ����� <^8�8 �r�l��� 4 � �X��� P �1� �X��4-� �X� P �&4 � ��4 ��pS�4p�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��@4 �?0 ��� p��P ��r�l�48��0P 48��*0.���r�l�48��$P 48��0@4�l48��                                            ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                4�l48��8�0 ��0�0��l4 �8�4�p�T�P ��8�4�h0 �8���P ��P��08�4�[8���p�Ip��0T��8���
8���
A P��4 �	�8��ۄ8��� 8 ���	B T��	8��΄	� �ր
��� ��� ��X��4� ��4	8��#�P�0�48 ��� ��� X��4 ���P�08���0�08���48��    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                ��8� �pT �
8��� t�� x��4 ��P4� �4 8 ��� X����8 ��8��4	8��_                                                                                                                                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0T4�l48��~8�0��l0�
0 �48��rP �B48��mP �8�4�h8���p�p��݀
P�
X�4� �
�P��'48��RP �"8�08�4�J�
8���0��
a 8���4 �	�	����� 8 ��A �	! 8���T��	8���08���48��&                                                                        