������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
 CAN'T OPEN FILE
                                                           0 ��� �<^8�8 �r�l��� 4 � �X��� P �.� �X��4-� �X� P �#4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��D4 �C0 ��� P ��4 �<                                                                                                              