������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: DEBUG FILE
 CAN'T CREATE FILE
 OUT OF SPACE
 BAD RECORD
 
?
@                                   0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ��� p��8Ȼ 48��:48��7                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0W�0Z8�4�l48��z4�l48��u0 ���	8�� 48��jP ��4��� 4 ��X ��pQ��P ��48��X�T �ӄ�	p�48��Op�48��Kp	48��G��0 ���4��� 4 ��X�40� �949� �4A� �34F� �0pp0���0E �J �Tp���H ��0���0��                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �P �A�	4�� �=8�8�� 48��t�	4��� 4 ��8�� 48��i0:48��g0�l48��b0 ��8�� 48��XP �P ��P ��T ��	�8��� 8 ��0���	P�	��48��>48��;                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �P �U�	4�� �Q8�8�� 48��t�	4	@ @ �T� ���� 8 ���8�� 48��b�8�� 48��\0:48��Z0�l48��U0 ��8�� 48��KP �P ��P ��	�8	@ @ �X� ��� 4 ������8 ��0���	P�	��48��*48��'                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �P �8�0�l�4	8��y48��t8��P �0�l�4	8��k�4���4@ �T� ��� T��8�� 4 ���	8�� 48��R48��O                                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0 �8 4��� 4��� X�����r�l�8�48��oP ��48��iP �0'�+0�l8 �
" 48��]P ��
0J4��� t��t���4@ �T� ��� T��4�� 0 ��X��0��\048��84 ��4�4�l48��1                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |4 ��4@ �T� ��� X �t��� 8 ���8�8�l48��jP �04 ���4���0� 0��04�� P��4��0 8 � P��4	��0 8 � P��4
��0 � P��0 ���0;T �	�
�P�
�0��\�54 ��4�4�l48��-                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8�0
48��}048��y�	8�� �0/48��q\�n|�� � � � 8�8�� �\�4� �p��4
� �PP04�W                                                                                                                                                                    