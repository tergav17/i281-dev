������������������������������������������������������������������������������������������������������������������������������HELLO, WORLD!
                                                                                                                 0 ��<^0�l0 48�8��x4 �w                                                                                                                                                                                                                                      