������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
 CAN'T OPEN FILE
                                                           0 ��� �<^8�8 �r�l��� 4 � �X��� P �.� �X��4-� �X� P �#4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��D4 �C0 ��� P ��0 �48��64 �74���                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8�� 48��{8�8�� 48��t�P ��48��n                                                                                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0��|0 ���0��P�� � ��r�l�8�8�48��lP �0�l0448��b4�l0 48��^P ��\�Y|�� � �'��P ���� 4 ��P��X �8
��0 T�8� ��P��8�48��6P �0 4���\��0 �\�)                                                                            