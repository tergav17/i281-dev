������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
                                                                                                               0 ��<^8�8�� 48��w�r�l��8 � 4 � �X��� P �� �X��� 4 �f                                                                                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 ����0 ���P ��0 �aX� ��`��`���m��0�T �h������ �< � ������0 �Y�������� �8 ������K                                                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8�48��}P �0 \�w                                                                                                                                                                                                                                          