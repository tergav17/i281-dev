������������������������������������������������������������������������������������������������������������������������������HELLO, WORLD!
                                                                                                                 4 � P ���J J J ����T����                                                                                                                                                                                                                                      