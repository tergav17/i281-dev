������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
  /FY 4Qh %6J^ (<                                    0 ����<^8�8 �r�l��� 4 � �X��� P �0� �X��4-� �X� P �%4 � ��4 ��pL�4T �0� �r�l����4 ����t�T���0 ��0�l0 8�48��B4 �A0 ���P ��0 �D0�N8һ 48��048��-4 �.4 ��� 48��%                                                                      ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
 UNEXPECTED CHAR IN NUMERIC
 UNDEFINED EXPRESSION
 UNEXPECTED TOKEN
 VALUE STACK OVERFLOW
                 8��G��
�r��� 4 ��4 � �48��t�
P��0:48��m�E��F�8�� �0:48��b0 48��^� p�@ P48��� �8 ���l48��N|8 �"0'48��04�8��0 4d8��0 4
8��00�"0 48��\�4�#�"����m �x�h ����< � �80�"X����P ��#�48��#�                              ������������������������������������������������������������������������������������������������������������������������������EXPRESSION STACK OVERFLOW
 VALUE STACK DEPLETION
 EXPRESSION STACK DEPLETION
 PARENTHESIS MISMATCH
 DIVIDE BY ZERO
        8�8�� 4	8��{8�� 48��v0 8�� 48��p0 �O�P8�8�� 4	8��f�;P �p
��pv48��]p48��Yp�48��U0�48��Q�DP �P�D��8�8�� 48��D48��A                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������OUT OF MEMORY
 LOCAL OUT OF RANGE
 FILE I/O ERROR
 TEXT SEGMENT FULL
 DATA SEGMENT FULL
 DATA IN BSS
                     04 D � 8��� 8��� 8��� 8 ��p��8�8�� 4	8��j�;p=�p��48��b8�� 48��]�Q�R�H���8 �0�� ���+8�� 48��M8�� 4	8��H8�� 48��CP �����Q�R����0�� 0 ����0 �Q�R��� ���;p
0�48��'48��$                                                                    ������������������������������������������������������������������������������������������������������������������������������UNKNOWN DIRECTIVE
 UNKNOWN DATA TYPE
 UNENCLOSED STRING
 VALUE OUT OF RANGE
                                                8�8�� 48��{�P ��4
� �0�48��p�DT �P08�� 48��g8�� 4	8��b�;p:�0�48��[�PP�P��OP�O48��Q                                                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������AOUT.SV CANNOT CREATE AOUT.SV
 ORG �TEXT �DATA �BSS �DEF �DEFL �BANK � BYTE WORD                                             8�8�� 4	8��{0 8�� �R�"8�� 4	8��q�"X �0��D4�h0 8��g08��d08��a8��_8��]�;p��0H8�� �1P �0��*�S�%�;p��0H8�� �$P �0���S8û 4	8��?�;p��0��8ͻ 48��5�Q�R�H���8 �0�� ��48��(48��%�4 � <��� � �	X �< ��PT���� \ �P��P� ��X ��0 < ����      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8�� 4	8��{�;P �Up
�Sp�8�� 4	8��o�;p"�p��
P
�4 ��8�� 48��`0��>8̻ 4	8��Y8�� 48��T�DT �P 0��.�IP ��Sp���"��0 �8Ż 48��=�"�8̻ 48��6�;p,�	8Ի 4	8��.�;p
�����;P �p
�0��48�� 48��                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8�� 48��{P 0��4��H�P 0��.�#�J�S8�8�� 48��hP 0��!��J�P 0���S�"�I8�� 48��W�J�"8�8�� 48��N�;P �p
�0��48��D48��A                                                                                                                              �	�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                |4
�8��@P�{�@8��x0��<0��C0��@|0 �?�=�A�B0�>�<P�<�� ��r�l�8	�8�48��]P �	�<�G0 �E�F0�48��P4�l0 48��LP ��\�G|�<�� �)�?�>P ���� 4 ��P�?�CX �8
�C�0 T�>8� ��=P��=4�l8	�48��"P �0 4�>��\��0 �C\�                                    �
�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                �<�G�BP�B�A�T�A�E�F�CP �l�=4
� �4��@�e�@4;� �3X �4 � �.40� �49� 4��,4a� �4z� �p 4_� �4A� �4Z� 4���@� �8 �@�>X �<4;� ��@�	4'� �4"� ��0�@�.8�� 4	8��1�;8 � �
8ڻ 4	8��(�
�C40� �49� �4a� �4z� �p 4_� �4A� �4Z� �X4� ����0 ��4��C�;\�  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0
�"0 ��0 � T �wt0�	4�"P� 89� �P�( � T �X����t9�T9�
0 ���
8tX�t��
8t�8t��0�48��N�"�
� P �J����"|�	�B ���PA �����
� P40� ��49� �4A� ��4F� ��xx0�"� �ӄF ��ԄT���                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                               |0 �:0.�90$�88�0 ��;p���P ��pB�p�0��O� �P�!� 8�� 48��`P �%�:�#8ɻ 48��Wp��	8�� 48��PP ��:�p��8��1�;�8��-�;p'�0�48��=p��H��903� 0���� ��T�9�p����80)� 0���;� ��T�8�0�48��8�8� 4	8���;�p���p���p���p��p���48��    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8p�<p�:8p��7p�5p��38pW�08p��-8p��*8p=�'p���84$� �0�48��^��t(�8�� 48��Vp�8�#p�p��"8�� 4	8��J�;�� 8�0�48��A��84$� �	���� �8» 48��348��048��-�84$� �8ջ 48��$�940� �0�48���������:\�                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0��88$� �ft�80��980� �_���!��� ������t�9�:P �L�8� p+���!A ��� �PA ��=p���!a ��� �pa ��0p��+���0 ��X �\ ���"� �� �\��� �\���!A ��� �PA ��!@ �!� �@ P� ��@ � ��48���9�������48��                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                p�p��O� P ��!P �0��P�8 < 0��@ ���	@ �P��Pp ��@ ��O �O �\�\| �J �J �X�Xx �!l � �x�h P �h ��!L �X� H ��P��p�ŀ8� p/�����48��,�9�������'48��#                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                p�� X 4��!� �& T �c�� ���� P���� �p��� X 4��!� �& T �L�@ ���@ P��@ �t��p���� 8@ �E �P�E x�����!8@ �E �P�E x����"pV��� 8@ �E P�E �Px�����!8@ �E P�E �Px����48���9�������                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                p���� 8@ �E �P�E �Px�����!8@ �E �P�E �Px����)p��!�� 4�f 8@ �E P�E �Px�����!4�f 8@ �E P�E �Px����p�0�48��8�9�������3                                                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��48��|�4<�"8�X� �"��� � �P �0 ��\x��8n \��� 8 ����0�c ��\n � P �\�|0 ���ـ P 8 ����"<��8 ���0��E�4 �"8<����� 4 ����!T �� T ��"�#�!t�!�� t� �4 � �!X��8��� \ ��4 ���T ��"�#0�\ ���� 0 ������                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �4<�Q8�X� �Q��� � �P �0 ��\x��8n \0 ���R��hn � P �&\�|0 ���߀ P 8 ����Q<�ׄN�q� �0�48��MT�Nt�Q��� ��0 8� � �X������8\4 ��|x�� �Q��� ��\	��                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                4) ��� T ���T�4 ����N�q� ��0�48��mT�Nt��� ) ��<�4 � � \��4 �����4t� 0 ���H���T�0 ���O                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 �L4 08��108��.|4�l0 8�48��rP �048��l4 �j0 �K\�e4 08��08���P �4�08��08���H0 �I0�J48��K��0 � P��0 ���A48��@48��=                                                                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |4�l0 8�48��{P 0�48��t�KP 48��o�M4@ �T� ��� X �t��� 0 ���8�� 8 ���LX�Lxt��� 0 ��" 4�l4	8��NP 0�48��G48��D                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8��J4@ �T� ��� X �t��� 0 ��" 4�l48��mP 0�48��f�4 ���J4���0� 0��04�� P��4 08��08��08���<�� ��r�l�48��DP 0�48��=�J�M0 �K\�8��0 � P��0 ���-                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |�DP �B�M�J� �8�8�� 48��s�IP ��H�T �p�P �0�48��e4@ @ �T� ���� 8 ������8 ����HP �0�48��M�I�t�X �0�48��C4��� 8 ��0��K�HP�H\�8                                                                                                          ������������������������������������������������������������������������������������������������������������������������������        NOOP  INPUTC INPUTD INPUTCF INPUTDF MOV  LOADI 0ADD @ADDI PSUB `SUBI pLOAD �LOADF �STORE �STOREF 	�   �I�IT �4�4�"@ �T� �H��� 0 ���IT �4�4�J@ �T� ��� 0 ���H�a                                                                                                                                                                                            ������������������������������������������������������������������������������������������������������������������������������        SHIFTL @SHIFTR 
�CMP �CACHE WRITE BANK  BRC �BRAE �BRNC �BRB �BRO �BRNO �BRN �BRNN �BRP �BRZ �BRE �   08�� �P �08���P �	08���P �0�48��n�S48��j���40 � � � �PT\ ��� ��\ �T� ��T� \ ��0 4 8 ���� �I|8��;p���P �� pA4� �	�"8˻ 4	8��7�"\�50�48��0                                                                                            ������������������������������������������������������������������������������������������������������������������������������        BRNZ �BRNE �BRA �BRBE �BRG �BRGE �BRL �BRLE �JUMPR �JUMP �NOR �NORI �                                       8�p�	�S�0 �8� 48��up�+8�� 48��n�S@ @ D �S�;p,�I8��>8����SD �S0 ��;p+�8��28�� 48��S�DT �P �0��4�S�8���p�8��҄S@ @ D �S�;p,�8��8ͻ 48��5�DT �P �0���S�8���48��'8� 4	8��"�;P �p
�0��48��48��                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�p��;p[�i8��^8�� 48��t�DT �P �0��`�S�8�� 48��f�;p]�Q�Fp��;p[�K8��@8�� 48��V�S@ @ D �S�;p+�8��1�S�0 �8���p�8���S@ @ D �S�;p,�(8��p�8��ڄS@ @ D �S�;p,�8���;p[�8��
8��ɄSD �S��48��8� 4	8���;P �p
�0��48��48��
                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�p�*�;p[�l8��a8�� 48��t�DT �P �0��c�;p]�[8��P�;p,�V8��K8�� 48��^�S@ @ D �8� 48��Tp��;p[�@8��58���SD �S0 ��;p+��8��)p�8��ۄS@ @ D �0 �8���p�8ջ 48��-�DT �P �0���S��H4�d �A �8���48��8� 4	8���;P �p
�0��48��
48��          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�p�8�� 48��y�S( @ @ D F �0 �8̻ 48��kp� 8���p�4��;p+�8��%8�� 48��Z�DT �P �0��'�S��H4�d �A �8���p�	8���P ���S�8���48��;8̻ 4	8��6�;P �p
�0��48��,48�                                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�p�9�;p[�`8��U8�� 48��tP �W�S@ @ D �S0 ��;p+�8��B8�� 48��a�DT �P �0��D�;p]�<8��1�;p,�78��,8���P �1�S�8� 48��Ep�(8��ɄS@ @ D �S0 ��;p+�8��8һ 48��0�DT �P �0���S�8���8� 4	8�� �;P �p
�0��48��48��                                  