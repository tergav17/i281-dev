������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: TEMPLT [-A] FILE1 FILE2 ...
 FAILED TO OPEN FILE
 FILE TOO LARGE
                                  0 ��� �<^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0 4�l48��G4 �F0 ��� p��r�l�48��:P 08��0 4��l48��0P �
��lPT�px� ��0N��48��                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�  48��~P ��48��y4 �x                                                                                                                                                                                                                                      