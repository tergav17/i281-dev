������������������������������������������������������������������������������������������������������������������������������?:*.*  FILES IN USE
  BLOCKS IN USE
  BLOCKS FREE
                                                                           0 ��<^48�8��{0 ����	0�l0 4
8��pP ��P���P��	�iA �	��P�hA ��	P�	��P�48��S�� ��08�� 48��G048��E�� �	�08Ȼ 48��9048��748��4�n� �o�08ٻ 48��(0'48��&4 �%                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8 �P �0'48��04�8��0 4d8��0 4
8��00�0 48��\�e����� �m �x�h �� ��< � �80�X����P ���F48���D                                                                                                                                  