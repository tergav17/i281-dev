������������������������������������������������������������������������������������������������������������������������������
?
%                                                                                                                          0 ��<^8���r�l��8 � 4 � �X��� P �� �	X��0 ��8�� 48��d<� 4 ��� p �X\4'� ��r����0 � �8�� 48��MP 48��I48��F4 �G                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 �08�4�l48��z4�l48��u0 ������0 ���4��� 4 ��P�0,� �*00� ��09� �+�P �0��
8	������D ����T��D ���x��
x0�B ���P���ˀp����0���" 4Q� 4 �+4F� 48��#�4��� 4 ��X ��48��                                            ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                4P� 48��}4R� 48��x4W� 48��s4A� 48��n4I� 48��i4D� 48��d4M� 48��_4L� 48��Z48��W48��T                                                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��48��|48��y48��v48��s48��p48��m�P �!��4��� X4 � �� � �<� 4 ��� p �X\4'� �4����0 � �48��I4 ��48��D48��A                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �p�Y�������� �P���� �K����8�8�� 4	8��fP �>� ���� 8 ��P �
�48��Z��T�� �� ���� �8 ��P � � �T�T��ހ�� ����� ��P���P��0
48��/048��+48��&48��#                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �P �58�8�� 48��xP �,�(�p�(��P �T ���8�8�� 4	8��cP �0�8�8�� 4	8��YP ��	�p���p��(��48��J48��G                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �p�%�������� ����� �����8�8�� 4	8��fP �
8�� 4	8��_P �48��Z48��W|8 �,0'48��04�8��0 4d8��0 4
8��00�,0 48��\�=�-�,�
���m �x�h ����
< � �80�,X�
���
P ��-�48��-�                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |�P �5�*�+��0
48�8��v048��r8�� 48��k\48��g|�P ����8 <��� �X ����0 ���A ���P���0 �����\48��E�P �8�8ǻ 48��;�48��9�P �48��148��.                                                                                        �	�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��4
8��|��0 �(0�)� �0�T �r���0 ��T ��( a ���t��P �T �
� ��(�)��� �0 ���ހ �T ��T��� P �T��x���0 ����B0 ��0��>                                                                                                                      �
�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                |�P �	0 4� �0�0 ��"� ���X� ���� \ ���� �P �8I ���	< ��� ��8 I ���< ���4�l48��P�0��� 0 ��T �7� �����8
�8ǻ 48��;P �+�� ��0 ���T8 0��� 0 ��� \ �����P�< ���� 0 ��TX\ ������ ��T �48��\�                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�0
48��~048��z48��w8��8�� 8��� �p.�T 8 ���^0 ���� T� ���� X 8 ����< � ���� P ��p�� 8��� 8��8 ��T\�� ��8 �0�X�����0 ��X ��T� �� ���� X ��X�0 ����
�8� 48��P ��8 ���
��p� �� ��0��0 ��4
8��	\�          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |���� �����p�0�� X \� �� P �0�������\ < ������x� ��(�)��� �8 ���8�8�� 48��Q���� ��(�)� �<M �8 I P �)��|��0 ������� ����� �	�P���P�������� � �
��� �� � <��PX��0 ���\�                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 �����0 ���P ��0 �aX� ��`��`��8f E �PE �@ P�*�+�b��T 0��]������ �< � �����0 ���P�P�0 ��+p�+��*p�*��� ������ ���� �0 ��� ���� �0 ����� �0 ��%�� ������ �8 �����+P�+��*P�*��                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8��	48��||8
�	0 �l08�48��sP �8�� 48��j0 � ��0�8�� 8�48��]\�\                                                                                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0�l0 8��48��{P �K0�4 �	�	tX �T���� 0 ���4 � �4�� �
�)4	� �X �04
� �!8 ��� � ���� 4 ��X ��T�P���
�����4 ���8Ȼ 48��:�
����T��4 P8� ���P������� ��� �<�� ��< ���0 4 ��\�                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�48��0 �l08�48��wP �V0�l�0�0 ����4G \ ��� �0 X ���� 4 ��P 4��0$ �
��\ �X<� < ���8�4	8��GP �&�P�0�� 8< �
T ���� 0 ��\��T ��t4
�ׄ� �T� �¨�����0 ��< M T��0 4 ���\�                                            