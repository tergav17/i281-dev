������������������������������������������������������������������������������������������������������������������������������
?
%                                                                                                                          0 ��<^8���r�l��8 � 4 � �X��� P �� �	X��0 ��8�� 48��c<� 4 ��� p �X\4'� ��r����0 � �8�� 48��LP 48��H48��E4 �F                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 ����0 ���P ��0 �aX� ��`��`���m��T 0��h������ �< � �����0 ���P�P�0 ���� ������ ���� �0 ��� ���� �0 ����� ���8�� ������ �8 ������*� �0�T �%��� �0 ��0�T �� �0 �                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8
�	0 �l08�48��xP �8�� 48��o0 � ��0�8�� 8�48��b\�a                                                                                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0�l0 8��48��zP �K0�4 �	�	tX �T���� 0 ���4 � �4�� �
�)4	� �X �04
� �!8 ��� � ���� 4 ��X ��T�P���
�����4 ���8Ȼ 48��9�
����T��4 P8� ���P������� ��� �<�� ��< ���0 4 ��\�                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 �08�4�l48��y4�l48��t0 ������0 ���4��� 4 ��P�0,� �*00� ��09� �+�P �0��
8	������D ����T��D ���x��
x0�B ���P���ˀp����0���0Q� 4 �+�4��� 4 ��P ��" 48��                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                4P� 48��|48��y48��v                                                                                                                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �p�Y�������� �P���� �K����8�8�� 48��eP �>� ���� 8 ��P �
�48��Y��T�� �� ���� �8 ��P � � �T�T��ހ�� ����� ��P���P��0
48��.048��*48��%48��"                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                ��� �0�T �{���0 ��T ��( a ���t��P �T �� ���� �0 ����� �T ��T��� P �T��x���0 ����M0 ��0��I                                                                                                                                              