������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: HDUMP FILE {START BLK} {END BLK}
 CAN'T OPEN FILE
 :                                                0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ���	0��
� P ��p��0̳ ��	�
� p��0ճ �
�
�	� �ۀ p��48��#0 �r��� t �t��t
��$ @ ��@ ��@ ��A ��A ��� t0A �X��4 ���4 �  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8��r�l�48��|P �0�l0=48��t8�0�l�	48��lP �/0�0 �4��	E 0�0 8�� 48��X�	@ �t�P8�� 48��M��t� �P�8�� 48��B0�l0O48��>48��948��6                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�0������ 8 ��8�� �'�T���p���0 48��k�p���8�0L48��a0 ��p�P���	�
� �P�	48��N|�� � � � 8�8�� �\�4� �p��4
� �PP04�848��2                                                                                                