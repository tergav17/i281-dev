������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
                                                                                                               0 ��<^8�8�� 48��w��r�l��8 � 4 � �X��� P �� �X��0 ���<� 4 ��� p �X\4� ��r����0 � �8�� 48��K4 �L                                                                                                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 �	�
��0 ���P ��0 �aX� ��`��`���m��	T 0��h�
����� �< � ����	�
0 ����������� ���� �0 ������� �0 ����C����	�
��� �8 ���	�
��5                                                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0 �l0��8�48��y��P ���8�� 48��n��0 ���0�8�� 48��b0�l0 � 48��]P � 0 \�W                                                                                                                                                                          