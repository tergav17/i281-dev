������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: SH FILE
 FILE NAME TOO LONG
                                                                        0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ��� p��48� ��r��� 8 ���s��� 8 ��PT| ��k�s��0�� �0 �����4 �"<^0�l0$48��                                            