������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: YMPLAY
                                                                                              0 ��� <^8�8 �r�l��� 4 � �X��� P �-� �X��4-� �X� P �"4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��F4 �E0 ��� P ��0 ��������4��4द4��0��0���0��0��48��%                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 ��	8�8��Q0 ��8��M8��4 ��� T��X0� ��0 ���P���P�������4��4द4��8��-0 ��0 4����� 4 ��8�� 48��HP �0����0������
��P��0 T8� ����0 ��8��0 ����P��4 �-��E ��E ���"                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                ( �t��	T�	0�t�xY�E�vt�xM�@�qt�x5�;�lt�x!�6�gt�30��0�t�|8�P �
�T�0 �	0
48��R048��N\��	�
T�	t�4 �	�
pE�	�pn��pd��p!�48��30��20 �0                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8��
�E @ �T�
���E @ �T����E @ �T����E @ �T���@ 4� �! ��@ @ � � P��8�
��������x��48��HP �0��    ��� ��0��0 ��0���0�\�40 \�1                                                                                            