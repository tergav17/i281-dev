������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
                                                                                                               0 ��<^8�8�� 48��w��r�l��8 � 4 � �X��� P �� �X��0 ���<� 4 ��� p �X\4� ��r����0 � �8�� 48��K4 �L                                                                                                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 �
���0 ���P ��0 �aX� ��`��`���m��
T 0��h���	��� �< � ����
�0 ��������	��� ���� �0 ������� �0 ����C����
���� �8 ���
���5                                                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0 �l08�48��zP �P8�� 48��q0 ���0�8�� 48��f�P�P �0 �0�l0 � 48��ZP �%04 ����� 0 ����� ����� 4 ��P��8Ļ 48��=��T��4 P8� ��� P�Հ��� ����4�� ��0 4 ��\�#                                                                  