������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
  /FY 4Qh                                                       0 ��� �<^8�8 �r�l��� 4 � �X��� P �0� �X��4-� �X� P �%4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��B4 �A0 ��� P ��0 �D0
�L48��24 �34 ���48��*                                                                                ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
 UNEXPECTED CHAR IN NUMERIC
 UNDEFINED EXPRESSION
 UNEXPECTED TOKEN
 VALUE STACK OVERFLOW
                 8��G��8�r��� 4 ��4 � �48��t�8P��0:48��m�E��F�8�� �0:48��b0 48��^�p�@ P48��� �8 ���l48��N|8 �0'48��04�8��0 4d8��0 4
8��00�0 48��\�4������m �x�h ����< � �80�X����P ���48���                              ������������������������������������������������������������������������������������������������������������������������������EXPRESSION STACK OVERFLOW
 VALUE STACK DEPLETION
 EXPRESSION STACK DEPLETION
 PARENTHESIS MISMATCH
 DIVIDE BY ZERO
        8�8�� 48��{0 �M8�8�� 48��r�/P �4p
��8�� 48��h8�� 48��c�/p=�0�48��\8�� 48��W8�� 48��RP �����O�P����0�� 0 �����0 �O�P��� ����0A�90 �:8�0A48��30=48��/8ڻ 48��(P �8� 48��!0?48��48��                                                ������������������������������������������������������������������������������������������������������������������������������OUT OF MEMORY
                                                                                                                 |4�8��4P�{�48��x0��00��50��4|0 �3�1�6�70�2�0P�0� � ��r�l�8�8�48��]P �	�0�G0 �E�F0�48��P4�l0 48��LP ��\�G|�0� � �'�3�2P ���� 4 ��P�3�5X �8
�5�0 T�28	� ��1P��18�48��$P �0 4�2��\��0 �5\�                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �0�G�7P�7�6�T�6�E�F�5P �l�=4
� �4��4�e�44;� �3X �4 � �.40� �49� 4��,4a� �4z� �p 4_� �4A� �4Z� 4���4� �8 �4�>X �<4;� ��4�	4'� �4"� ��0�4�.8�� 48��1�/89� �88ڻ 48��(�8�540� �49� �4a� �4z� �p 4_� �4A� �4Z� �X4C� ����0 ��4��5�/\�  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0
�0 ��09� T �wt0�	4�P� 89� �P�( � T �X����t9�T9�80 ���88tX�t��
8t�8t��0�48��N��8� P �J����|�	�B ���PA �����8� P40� ��49� �4A� ��4F� ��xx0�� �ӄF ��ԄT���                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0 �.0"�-0�,8��/p���;P �	�:pF�p��0 ���8�� 48��ep��	8�� 48��^P ��.�p��0 ��H��-0'� 0���� ��T�-�p����,0� 0���/� ��T�,�0�48��58�8Ի 48��.�/�p���p���p���p���48��!                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8p�<p�:8p��7p�5p��38pW�08p��-8p��*8p=�'p���,4� �0�48��^��t(�8�� 4	8��Vp�,�#p�p��"8�� 48��J�/�� 8�0�48��A��,4� �	���� �8» 4	8��348��048��-�,4� �8ջ 4	8��$�-4$� �0�48���������.\�                                      �	�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                0��,8� �ft�,0��-8$� �_������������t�-�.P �L�,� p+���A ����PA ��=p���a ����pa ��0p��+���0 ��X �\ ���"� �� �\��� �\���A ����PA ��@ ���@ P���@ ���4
8���-�������48��                                    �
�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                p�p��O�P ��P �0��P�8 < 0��@ ���	@ �P��Pp ��@ ��O �O �\�\| �J �J �X�Xx �l ��x�h P �h ��L �X�H ��P��p�ŀ,� p/�����48��,�-�������'48��#                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                p��X 4��� �& T �c�� ���� P���� �p���X 4��� �& T �L�@ ���@ P��@ �t��p����8@ �E �P�E x�����8@ �E �P�E x����"pV���8@ �E P�E �Px�����8@ �E P�E �Px����48���-�������                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                p����8@ �E �P�E �Px�����8@ �E �P�E �Px����)p��!��4�f 8@ �E P�E �Px�����4�f 8@ �E P�E �Px����p�0�48��8�-�������3                                                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48���4	<�8�X�9���� � �P �0 ��\x��8n \��� 8 ����0�c ��_n � P �\�|0 ���ـ P 8 ����<��8 ���0��H                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �4	<�O8�X�9�O��� � �P �0 ��\x��8n \0 ���P��hn � P �&\�|0 ���߀ P 8 ����O<�ׄL�q� �0�48��MT�Lt�O��� ��0 8� � �X������8\4 ��|x��9�O��� ��\	��                                                                                          