������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: DEBUG FILE
 CAN'T OPEN FILE
 CAN'T CREATE FILE
 
?
*                                             0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ��� p��48��<��                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0M�0P8�4�l48��z4�l48��u0 ���	8�� 48��jP ��4���4 ��X ��pQ48��\p�����0 ���4��� 4 ��X�40� �L49� �4A� �F4F� �Cpp0���0E �J �Tp���H ��0���0��-                                                                                    