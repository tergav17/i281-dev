������������������������������������������������������������������������������������������������������������������������������NO ARGUMENT
 CAN'T OPEN FILE
                                                                                                 0 ��<^8��r�l��8 � 4 � �X��� P �� �
X��0 ��0�l0 48��f0 ��" 48��`P �0�l048��X0�l0 � 48��QP �0 4����� P �4 ��48��B��P��0 T8� �� P��4 �5                                                                                                