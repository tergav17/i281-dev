������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: CAT FILE1 FILE2 ...
 CAN'T OPEN FILE
 PRINTER NOT READY
                                           0 ��� �<^8�8 ��r�l��� 4 � �X��� P �.� �X��4-� �X� P �#4 � ��4 ��pP�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��C4 �B0 ��� P ��48��7                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8��P �0 �48��zP �	�P ��0�l0B48��o�r�l��48��hP �0�l0048��`0�l0 �48��YP �0 4����� P �4 ���T �48��G48��D��P��0 T8� ��P��4 ���P�� � ��4 �/                                                                                    