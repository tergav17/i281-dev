������������������������������������������������������������������������������������������������������������������������������
?
%                                                                                                                          0 ��<^8���r�l��8 � 4 � �X��� P �� �	X��0 ��8�� 48��d<� 4 ��� p �X\4'� ��r����0 � �8�� 48��MP 48��I48��F4 �G                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 ����0 ���P ��0 �aX� ��`��`���n��T 0��i������ �< � �����0 ���P�P�0 ���� ������ ���� �0 ��� ���� �0 ����� ���9�� ������ �8 ������+� �0�T �&��� �0 ��0�T �� �0 �                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8
�	0 �l08�48��yP �8�� 48��p0 � ��0�8�� 8�48��c\�b                                                                                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0�l0 8��48��{P �K0�4 �	�	tX �T���� 0 ���4 � �4�� �
�)4	� �X �04
� �!8 ��� � ���� 4 ��X ��T�P���
�����4 ���8Ȼ 48��:�
����T��4 P8� ���P������� ��� �<�� ��< ���0 4 ��\�                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 �08�4�l48��z4�l48��u0 ������0 ���4��� 4 ��P�0,� �*00� ��09� �+�P �0��
8	������D ����T��D ���x��
x0�B ���P���ˀp����0���" 4Q� 4 �+4F� 48��#�4��� 4 ��X ��48��                                            ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                4P� 48��}48��z48��w                                                                                                                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �P �48��|48��y48��v                                                                                                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �p�Y�������� �P���� �K����8�8�� 4	8��fP �>� ���� 8 ��P �
�48��Z��T�� �� ���� �8 ��P � � �T�T��ހ�� ����� ��P���P��0
48��/048��+48��&48��#                                                                  �	�����������������������������������������������������������������������������������������������������������������������������                                                                                                                                ��� �0�T �|���0 ��T ��( a ���t��P �T �� ���� �0 ����� �T ��T��� P �T��x���0 ����N0 ��0��J                                                                                                                                              