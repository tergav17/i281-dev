������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: TEMPLT [-A] FILE1 FILE2 ...
 FAILED TO OPEN FILE
 FILE TOO LARGE
                                  0 ��� �<^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0 4�l48��G4 �F0 ��� p��r�l�48��:P 08��0 4��l48��0P �
��lPT�px� ��0N��48��                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�8�� 48��{8�� 48��v8�� 48��q48��pP ��48��k4 �j                                                                                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������

	                                                                                   �������                                                                                                                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������]��<�s�k��N��O�u5���W'�ϧ�];��Ŭ�}hS@.����ʾ������xqke_ZUPLGC@<9520-*(&$"                                                                                                                                                                                                                                                                                                 