������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
                                                                                                               0 ��<^8�8�� 48��w�r�l��8 � 4 � �X��� P �� �X��0 ����<	� 4 ��� p �X\4� ��r����0 � �4 �Q                                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 ����0 ���P ��0 �aX� ��`��`���m��0�T �h������ �< � ������0 �Y�������� �8 ������K                                                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0 �l0`8�48��zP �0 \�t                                                                                                                                                                                                                                    