������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 ��<^48�8��{0�l04
8��u048��q�j4���4 ��048��g0�0 � �`48��_� �P� ���p�0.48��S0�0��0 48��K8�� 48��D0 48��B48��?P ��4 �<                                                                                                                ������������������������������������������������������������������������������������������������������������������������������
 UA NAME   EX SIZE
 0:  *.* NO FILES
                                                                                       � |8 �P �0'48��04�8��0 4d8��
0 4
8��0 48��\�f����h�im �x�h ��h�i�< � �80�X���48���K                                                                                                                                                