������������������������������������������������������������������������������������������������������������������������������NO ARGUMENT
 CAN'T REMOVE FILE
                                                                                               0 ��<^0�� 8��r��8 � 4 � �X��� P �� �
X��0 ��0�l0 48��e0 ����r�l�48��\P �48��WP �	� P �	0�l048��L0 � ��4 �H                                                                                                                                      