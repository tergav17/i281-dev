������������������������������������������������������������������������������������������������������������������������������HELLO, WORLD!
                                                                                                                 0 ��<^0�l0 48�8��y4 �x                                                                                                                                                                                                                                      