������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
                                                                                                               0 ��<^8�8�� 48��w��r�l��8 � 4 � �X��� P �� �X��0 ���<� 4 ��� p �X\4� ��r����0 � �8�� 48��K4 �L                                                                                                                                                ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8�q0 ����0 ���P ��0 �aX� ��`��`���m��T 0��h��
���� �< � �����0 ���P�P�0 �����	�
���� ���� �0 ����	��� �0 ����<���	����� �8 ������.                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8
�0 �l08�48��xP �8�� 48��o0 ���0�	8�� 8�48��b\�a                                                                                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0�l0 8�� 48��zP �I0�4 ��tX �T���� 0 ���4 � �4�� ��'4	� �	X �.4
� ��T�8 ��� ����� 4 ��P����	����4 ���8ƻ 48��;����T��4 P8� �À P������ ����4�� ��0 4 ��\�                                                          