������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: DEBUG FILE
 CAN'T CREATE FILE
 OUT OF SPACE
 BAD RECORD
 
?
*                                   0 ��� <^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��H4 �G0 ��� p��48��<��                                                                                                                  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0W�0Z8�4�l48��z4�l48��u0 ���	8�� 48��jP ��4���4 ��X ��pQ48��\��0 ���4��� 4 ��X�40� �N49� �4A� �H4F� �Epp0���0E �J �Tp���H ��0���0��/                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 8 4��� 4��� X�����r�l�8�48��qP �48��lP �0'�0�l0 �
48��aP ��
0J4��� t��t���4J �T� ��� 4�4�l48��F                                                                                                                                    