������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: XMODEM [-ST] FILE
 CAN'T OPEN FILE
 CAN'T CREATE FILE
 TRANSFER FAILED
                           0 ����� <^8�8 �r�l��� 4 � �X��� P �1� �X��4-� �X� P �&4 � ��4 ��pS�4p�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��@4 �?0 ��� p��P 48��2��                                                                                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �r�l�8�48��|P �0@4�l48��t0 �0��l4 �	8�4�j�	T�P ��8�4�b0 �	8���P ��	P��08�4�U8���p�?p��0T��8���8���A P��4 �
�8��ۄ8��� 8 ���
B T��
8��΄
� ���4� ��4	8��'�P�0�48 ��� ��� X��4 ���P�08���0�08���48��            ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                ��8� �pT �
4 8��� p�� x����P4� �4 8 ��� X����8 ��8��4	8��_                                                                                                                                                                                      