������������������������������������������������������������������������������������������������������������������������������NO ARGUMENT
 INVALID USER AREA
                                                                                               0 ��<^8��r�l��8 � 4 � �X��� P �� �
X��0 ��0�l0 48��f40� �49� ��4:� �	�4 � �� 4 ���k�0 ��0�l048��K4 �J                                                                                                                                          