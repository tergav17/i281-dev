������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
                                                                          0 ��� �<^8�8 �r�l��� 4 � �X��� P �0� �X��4-� �X� P �%4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��B4 �A0 ��� P ��0 �048��44 �54 ���448��,                                                                                    ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
 UNEXPECTED CHAR IN NUMERIC
                                                                                  8�8�� 48��{8�8�� 48��t�P �p���8�� 48��j��48��f                                                                                                                                                                                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                8��3��$�r��� 4 ��4 � �48��t�$P��0:48��m�1��2�8�� �0:48��b0 48��^�4p�@ P48��� �8 ���l48��N|8 �0'48��04�8��0 4d8��0 4
8��00�0 48��\�4������m �x�h ����< � �80�X����P ���48���                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0��0��!0�� |0 ���"�#0��P�� � ��r�l�8�8�48��dP �	��30 �1�20�48��W4�l0 48��SP ��\�N|�� � �'��P ���� 4 ��P��!X �8
�!�0 T�8� ��P��8�48��+P �0 4���\��0 �!\�                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |8�� P�� ��3�#P�#�"�T�"�1�2�!P �f�:4
� �4�� �_� 4;� �0X �4 � �+40� �49� 4��)4a� �4z� �p 4A� �4Z� 4��� � �8 � �;X �94;� �� �	4'� �4"� ��-� �+8�� 48��-�8%� �$8޻ 48��$�$�!40� �49� �4a� �4z� �p 4A� �4Z� �X4/� ����0 ��4��!�\�������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0
�0 ��0%� T �zt0�	4�P� 89� �P�( � T �X����t9�T9�$0 ���$8tX�t��
8t�8t��0�48��Q��$��N                                                                                                                                                      