������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: MLOAD FILE1 FILE2 ...
 CANNOT OPEN FILE
                                                            0 ��� <^8�8 �r�l��� 4 � �X��� P �-� �X��4-� �X� P �"4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��F4 �E0 ��� P ��0 ��48��7                                                                                                          ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                0 ��r�l�8�48��zP �0�l0248��r4 �q0�l0 �48��iP �'������4��4द4��8��"00��8��8��4 � ��T��X0� ��0 ���P���P��P�Ӏ� P� ��4 �:��E ��E ���/                                                                                              