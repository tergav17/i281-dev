������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: RM FILE
 CAN'T REMOVE FILE
                                                                         0 ��� 0��<^8�8 �r�l��� 4 � �X��� P �+� �X��4-� �X� P � 4 � ��4 ��T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 48��F4 �E0 ��� p��r�l�48��9P �48��4P �	�P �	0�l0$48��)0 ���4 �%                                                                