������������������������������������������������������������������������������������������������������������������������������INVALID ARGUMENTS
USAGE: AS [-L] FILE1 FILE2 ...
  /FY                                                                 0 ��� �<^8�8 �r�l��� 4 � �X��� P �0� �X��4-� �X� P �%4 � ��4 ��pL�4T �0� �r�l����4 ��� �t�T� ��0 ��0�l0 8�48��B4 �A0 ��� P ��0 �F48��44 �54 ���J48��,                                                                                    ������������������������������������������������������������������������������������������������������������������������������CAN'T OPEN FILE
 UNEXPECTED CHAR IN NUMERIC
 UNDEFINED EXPRESSION
 UNEXPECTED TOKEN
 VALUE STACK OVERFLOW
                 8�8�� 48��{8�8�� 48��t�1��P ���48��l                                                                                                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������EXPRESSION STACK OVERFLOW
                                                                                                     8��I��:�r��� 4 ��4 � �48��t�:P��0:48��m�G��H�8�� �0:48��b0 48��^�Jp�@ P48��� �8 ���l48��N|8 �0'48��04�8��0 4d8��0 4
8��00�0 48��\�4������m �x�h ����< � �80�X����P ���48���                              ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |4�8��6P�{�68��x0��20��70��6|0 �5�3�8�90�4�2P�2� � ��r�l�8�8�48��]P �	�2�I0 �G�H0�48��P4�l0 48��LP ��\�G|�2� � �'�5�4P ���� 4 ��P�5�7X �8
�7�0 T�48� ��3P��38�48��$P �0 4�4��\��0 �7\�                                        ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                �2�I�9P�9�8�T�8�G�H�7P �l�=4
� �4��6�e�64;� �3X �4 � �.40� �49� 4��,4a� �4z� �p 4_� �4A� �4Z� 4���6� �8 �6�>X �<4;� ��6�	4'� �4"� ��0�6�.8�� 48��1�18;� �:8ڻ 48��(�:�740� �49� �4a� �4z� �p 4_� �4A� �4Z� �X4E� ����0 ��4��7�1\�  ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                48��0
�0 ��0;� T �wt0�	4�P� 89� �P�( � T �X����t9�T9�:0 ���:8tX�t��
8t�8t��0�48��N��:� P �J����|�	�B ���PA �����:� P40� ��49� �4A� ��4F� ��xx0�� �ӄF ��ԄT���                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                |0#�00�/8��1p���=P �	�<pF�p��0 ���8�� 48��gp��0 ���p��0 ���00)� 0���� ��T�0�p��
�/0#� 0���1� T�0�0�48��@8�8ɻ 48��9�1p���p���p���p���48��-                                                                                      ������������������������������������������������������������������������������������������������������������������������������                                                                                                                                p�p�p��p�p��pV�	p��p��p9�p�� p                                                                                                                                                                                                                      